[translated]
module main

fn show () {
  if x := 5 > 3 {
    println((x).str())
}

}
fn main () {
  show()
}
