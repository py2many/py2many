@[translated]
module main

fn show() {
	x := 5
	if x > 3 {
		println(x.str())
	}
}

fn main() {
	show()
}
