module main

fn main() {
	println('Hello world!')
	println('Hello world!')
}
