@[translated]
module main

import math

fn main_func() {
	a := int(math.pow(2, 4))
	println(a.str())
}

fn main() {
	main_func()
}
