@[translated]
module main

fn main_func() {
	a := 2 ^ 4
	println(a.str())
}

fn main() {
	main_func()
}
