[translated]
module main

fn baz1() string {
	return 'foo'
}
