[translated]
module main

fn bar1() int {
	return 0
}
