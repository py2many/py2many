module main

fn main() {
	println('OK')
	exit(1)
}
